library ieee;
use ieee.std_logic_1164.all;

entity mips_control is
    port(   opcode              : in std_logic_vector(5 downto 0);
            funct               : in std_logic_vector(5 downto 0);
            RegDst, ALUSrc      : out std_logic;
            Jump, Jal, Jr       : out std_logic;
            Beq, Bne            : out std_logic;
            MemRead, MemWrite   : out std_logic;
            RegWrite, MemtoReg  : out std_logic;
            ALUControl          : out std_logic_vector(3 downto 0) );
end mips_control;

architecture arch of mips_control is begin
    process(opcode, funct) is begin
        case (opcode) is
            when "000000" =>
                case (funct) is
                    -- R TYPES
                    when "10" & X"0" => -- add (0x20)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "0010";
                    when "10" & X"1" => -- addu (0x21)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "0010";
                    when "10" & X"4" => -- and (0x24)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "0000";
                    when "00" & X"8" => -- jr (0x08)
                        RegDst      <=  '-';
                        ALUSrc      <=  '-';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '1';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '0';
                        MemtoReg    <=  '-';
                        ALUControl  <=  "----";
                    when "10" & X"7" => -- nor (0x27)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "1100";
                    when "10" & X"5" => -- or (0x25)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "0001";
                    when "10" & X"A" => -- slt (0x2a)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "0111";
                    when "00" & X"0" => -- sll (0x00)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "1000";
                    when "00" & X"2" => -- srl (0x02)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "1001";
                    when "00" & X"4" => -- sllv (0x04)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "1010";
                    when "00" & X"6" => -- srlv (0x06)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "1011";
                    when "10" & X"2" => -- sub (0x22)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "0110";
                    when "10" & X"3" => -- subu (0x23)
                        RegDst      <=  '1';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '1';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "0110";
                    when others =>
                        RegDst      <=  '0';
                        ALUSrc      <=  '0';
                        Jump        <=  '0';
                        Jal         <=  '0';
                        Jr          <=  '0';
                        Beq         <=  '0';
                        Bne         <=  '0';
                        MemRead     <=  '0';
                        MemWrite    <=  '0';
                        RegWrite    <=  '0';
                        MemtoReg    <=  '0';
                        ALUControl  <=  "0000";
                end case; 
            when "00" & X"8" => -- addi
                RegDst      <=  '0';
                ALUSrc      <=  '1';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '1';
                MemtoReg    <=  '0';
                ALUControl  <=  "0010";
            when "00" & X"9" => -- addiu
                RegDst      <=  '1';
                ALUSrc      <=  '0';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '1';
                MemtoReg    <=  '0';
                ALUControl  <=  "0010";
            when "00" & X"C" => -- andi
                RegDst      <=  '1';
                ALUSrc      <=  '0';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '1';
                MemtoReg    <=  '0';
                ALUControl  <=  "0000";
            when "00" & X"4" => -- beq
                RegDst      <=  '-';
                ALUSrc      <=  '0';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '1';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '0';
                MemtoReg    <=  '-';
                ALUControl  <=  "0110";
            when "00" & X"5" => -- bne
                RegDst      <=  '-';
                ALUSrc      <=  '0';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '1';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '0';
                MemtoReg    <=  '-';
                ALUControl  <=  "0110";
            when "00" & X"2" => -- j
                RegDst      <=  '-';
                ALUSrc      <=  '-';
                Jump        <=  '1';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '0';
                MemtoReg    <=  '-';
                ALUControl  <=  "----";
            when "00" & X"3" => -- jal 
                RegDst      <=  '-';
                ALUSrc      <=  '-';
                Jump        <=  '1';
                Jal         <=  '1';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '1';
                MemtoReg    <=  '-';
                ALUControl  <=  "----";
            when "00" & X"F" => -- lui
                RegDst      <=  '0';
                ALUSrc      <=  '1';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '1';
                MemtoReg    <=  '0';
                ALUControl  <=  "1101";
            when "10" & X"3" => -- lw (0x23)
                RegDst      <=  '0';
                ALUSrc      <=  '1';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '1';
                MemWrite    <=  '0';
                RegWrite    <=  '1';
                MemtoReg    <=  '1';
                ALUControl  <=  "0010";
            when "00" & X"D" => -- ori
                RegDst      <=  '0';
                ALUSrc      <=  '1';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '1';
                MemtoReg    <=  '0';
                ALUControl  <=  "0001";
            when "00" & X"A" => -- slti
                RegDst      <=  '0';
                ALUSrc      <=  '1';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '1';
                MemtoReg    <=  '0';
                ALUControl  <=  "0111";
            when "10" & X"B" => -- sw (0x2b)
                RegDst      <=  '-';
                ALUSrc      <=  '1';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '1';
                RegWrite    <=  '0';
                MemtoReg    <=  '-';
                ALUControl  <=  "0010";
            when others =>
                RegDst      <=  '0';
                ALUSrc      <=  '0';
                Jump        <=  '0';
                Jal         <=  '0';
                Jr          <=  '0';
                Beq         <=  '0';
                Bne         <=  '0';
                MemRead     <=  '0';
                MemWrite    <=  '0';
                RegWrite    <=  '0';
                MemtoReg    <=  '0';
                ALUControl  <=  "0000";
        end case;
    end process;
end arch;